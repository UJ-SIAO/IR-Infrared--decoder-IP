`timescale 1ns/1ns

module edge_detect_tb;

parameter BIT_PERIOD      = 8680; // (1/115200)*1000000000

reg clk_50M;
reg rst_n;
reg data_in;
wire pos_edge;
wire neg_edge;

integer ii;

edge_detect u1 (
    clk_50M,
    rst_n,
    data_in,
    pos_edge,
    neg_edge
    );

always
  #10 clk_50M = ~clk_50M;
  
initial
  begin
  rst_n = 0;  
  data_in = 1;
  clk_50M = 0 ;
  #30 rst_n = 1;
  
  #133 data_in = 0;
  #211 data_in = 1;
  
  #319 data_in = 0;
  #113 data_in = 1;
  
  #100
      
  $stop;
  end
  

initial
  begin
  $monitor("time=%3d rst_n=%d data_in=%d pos_edge=%d neg_edge=%d",$time,rst_n,data_in,pos_edge,neg_edge);
  end
  
endmodule